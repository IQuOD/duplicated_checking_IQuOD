netcdf sample {
dimensions:
    depth = unlimited;   // Or specify an upper limit if known

variables:
    float z(depth);              // Depth below sea level in meters
        z:units = "meters";
        z:long_name = "depth_below_sea_level";
        z:valid_range = 0.0f, 11000.0f;
        z:positive = "down"	
        z:_FillValue = NaN;

    float Temperature(depth);    // Temperature in degrees Celsius
        Temperature:units = "degrees_Celsius";
        Temperature:long_name = "sea_water_temperature";
        Temperature:valid_range = -2.0f, 50.0f;
        Temperature:_FillValue = NaN;

    float Salinity(depth);       // Salinity in PSU (Practical Salinity Units)
        Salinity:units = "PSU";
        Salinity:long_name = "sea_water_salinity";
        Salinity:valid_range = 0.0f, 45.0f;
        Salinity:_FillValue = NaN;

    float Oxygen(depth);                // Oxygen concentration in mL/L
        Oxygen:units = "Micromole per kilogram (µmol/kg)";
        Oxygen:long_name = "Sea water dissolved oxygen";
        Oxygen:valid_range = 0.0f, 1000.0f;
        Oxygen:_FillValue = NaN;

    float Chlorophyll(depth);           // Chlorophyll concentration in mg/m^3
        Chlorophyll:units = "Microgram per liter (µg l-1)";
        Chlorophyll:long_name = "Chlorophyll";
        Chlorophyll:valid_range = 0.0f, 50.0f;
        Chlorophyll:_FillValue = NaN;

    int wod_unique_cast;         // WOD unique cast identifier
        wod_unique_cast:long_name = "WOD Unique Cast Identifier";
        wod_unique_cast:valid_range = unlimited; 
        wod_unique_cast:_FillValue = -9999;

    float lat;                   // Latitude in decimal degrees
        lat:units = "degrees_north";
        lat:long_name = "Latitude";
        lat:valid_range = -90.0f, 90.0f;
        lat:_FillValue =NaN;

    float lon;                   // Longitude in decimal degrees
        lon:units = "degrees_east";
        lon:long_name = "Longitude";
        lon:valid_range = -180.0f, 180.0f;
        lon:_FillValue = NaN;

    double time;                 // Time of data collection in seconds since 1970-01-01 00:00:00 UTC
        time:units = days since 1770-01-01 00:00:00 UTC";
        time:long_name = "Time";
        time:valid_range = unlimited; 
        time:_FillValue = NaN;

    string country;              // Country name where data was collected
        country:long_name = "Country";
        country:comment = "https://www.ncei.noaa.gov/access/world-ocean-database/CODES/country-list.html"
        country:_FillValue = "";

    string Temperature_Instrument;  // Device used for temperature measurement
        Temperature_Instrument:long_name = "Temperature Instrument";
        Temperature_Instrument:comment = "https://www.ncei.noaa.gov/access/world-ocean-database/CODES/s_29_probe_type.html"
        Temperature_Instrument:_FillValue = "";

    string need_z_fix;           // Instruction for fixing depths
        need_z_fix:long_name = "Need Z Fix for XBT bias correction";
        need_z_fix:comment = "https://www.ncei.noaa.gov/access/world-ocean-database/CODES/s_54_needs_depth_fix.html"
        need_z_fix:_FillValue = "";

    string Recorder;             // Device which recorded measurement
        Recorder:long_name = "Recorder";
        Recorder:comment = "https://www.ncei.noaa.gov/access/world-ocean-database/CODES/s_32_recorder.html"
        Recorder:_FillValue = "";

    float GMT_time;              // GMT time of data collection
        GMT_time:units = "hours";
        GMT_time:long_name = "GMT Time";
        GMT_time:valid_range = 0.0f, 24.0f;
        GMT_time:_FillValue = NaN;

    int WMO_ID;                  // WMO identification code
        WMO_ID:long_name = "WMO_identification_code";
        WMO_ID:valid_range = 0, 999999;
        WMO_ID:_FillValue = NaN;

    string dbase_orig;           // Database from which data were extracted
        dbase_orig:long_name = "Database of Origin";
        dbase_orig:_FillValue = "";

    string Project;              // Name of the project
        Project:long_name = "Project";
        Project:comment = "name or acronym of project under which data were measured"
        Project:_FillValue = "";

    string platform;             // Name of platform from which measurements were taken
        platform:long_name = "Platform";
        platform:comment = "https://www.ncei.noaa.gov/access/world-ocean-database/CODES/s_3_platform.html"
        platform:_FillValue = "";

    string Ocean_Vehicle;        // Ocean vehicle used for data collection
        Ocean_Vehicle:long_name = "Ocean Vehicle";
        Ocean_Vehicle:comment = "https://www.ncei.noaa.gov/access/world-ocean-database/CODES/s_74_ocean_vehicle.html"
        Ocean_Vehicle:_FillValue = "";

    int Access_no;               // NODC accession number (used to find original data at NODC)
        Access_no:long_name = "NODC_accession_number";
        Access_no:comment = "https://www.ncei.noaa.gov/access/world-ocean-database/CODES/s_1_accession.html"
        Access_no:_FillValue =NaN;

    string Institute;            // Name of the institute which collected data
        Institute:long_name = "Institute";
        Institute:_FillValue = "";

    string WOD_cruise_identifier;  // Two byte country code + WOD cruise number (unique to country code)
        WOD_cruise_identifier:long_name = "WOD Cruise Identifier";
        WOD_cruise_identifier:comment = "Two byte country code + WOD cruise number (unique to country code)"
        WOD_cruise_identifier:_FillValue = "";

    string dataset;              // WOD dataset identifier
        dataset:long_name = "WOD_dataset";
        dataset:comment = "https://www.ncei.noaa.gov/access/world-ocean-database/CODES/wod-datasets.html"
        dataset:_FillValue = "";

// Note: If a specific data field does not have information, please set it to its default value.

data example:

z = 100.0, 200.0, 300.0;
Temperature = 15.5, 16.0, 16.5;
Salinity = 35.0, 35.1, 35.2;
Oxygen = 5.5, 5.6, 4.6
Chlorophyll = 2.3, 2.4, 3.5;
wod_unique_cast = 12345678;
lat = -27.4698;
lon = 153.0251;
time = 92710.26;
country = "Australia";
Temperature_Instrument = "CTD: TYPE UNKNOWN";
need_z_fix = "";
Recorder = "RecorderModel123";
GMT_time = 14.58;
WMO_ID = 3901273;
dbase_orig = "US GODAE server (Argo)";
Project = "U.S. ARGO PROJECT";
platform = "Research Vessel";
Ocean_Vehicle = "SOLO-II (MRV Systems)";
Access_no = 42682;
Institute = "CSIRO";
WOD_cruise_identifier = "US038425";
dataset = "profiling float";
}
